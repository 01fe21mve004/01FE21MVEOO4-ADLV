Driver class
Class driver;
no_transactions;
virtual int_vif;
mailbox transaction gen2_driv;
int f (“mailbox_virtual _vif count/n”);
this .gen2_driv=gen2_driv;
this. mailbox = mailbox;
endfunction
task rset
